module Cnt_4b(

	);

