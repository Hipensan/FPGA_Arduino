module IMEM(
	input [15:0] i_PC,
	output [15:0] o_Inst
	);

reg [15:0] r_Inst[0:15];

initial
begin
	r_Inst[0] = 16'b1000000110000000;  
	r_Inst[1] = 16'b0010110010110010;  
	r_Inst[2] = 16'b1101110001100111;  
	r_Inst[3] = 16'b1101110111011001;  
	r_Inst[4] = 16'b1111110110110001;  
	r_Inst[5] = 16'b1100000001111011; 
	r_Inst[6] = 16'b0000000000000000;  
	r_Inst[7] = 16'b0000000000000000;  
	r_Inst[8] = 16'b0000000000000000;  
	r_Inst[9] = 16'b0000000000000000;  
	r_Inst[10] = 16'b0000000000000000;  
	r_Inst[11] = 16'b0000000000000000;  
	r_Inst[12] = 16'b0000000000000000;  
	r_Inst[13] = 16'b0000000000000000;  
	r_Inst[14] = 16'b0000000000000000;  
	r_Inst[15] = 16'b0000000000000000; 
end

assign o_Inst = r_Inst[i_PC >> 1];
endmodule